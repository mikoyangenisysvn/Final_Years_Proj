// ====================== TOP MODULE ======================
module pwm_top #(
    parameter WIDTH = 16
)(
    input  wire                 clk,
    input  wire                 rst_n,

    // Giao diện ghi/đọc register
    input  wire                 wr_en,
    input  wire                 rd_en,
    input  wire [3:0]           addr,
    input  wire [WIDTH-1:0]     wr_data,
    output wire [WIDTH-1:0]     rd_data,

    output wire                 PWM_OUT
);

    // ------------------- Wire kết nối -------------------
    wire              en;
    wire              mode;
    wire [WIDTH-1:0]  period;
    wire [WIDTH-1:0]  duty;
    wire [WIDTH-1:0]  prescaler_div;

    wire              slow_clk;
    wire [WIDTH-1:0]  cnt_val;

    // ------------------- Register Block -------------------
    pwm_register #(.WIDTH(WIDTH)) u_reg (
        .clk          (clk),
        .rst_n        (rst_n),
        .wr_en        (wr_en),
        .rd_en        (rd_en),
        .addr         (addr),
        .wr_data      (wr_data),
        .rd_data      (rd_data),

        .en           (en),
        .mode         (mode),
        .period       (period),
        .duty         (duty),
        .prescaler_div(prescaler_div)
    );

    // ------------------- Prescaler -------------------
    prescaler u_prescaler (
        .clk       (clk),
        .rst_n     (rst_n),
        .div       (prescaler_div[15:0]),   // chỉ dùng 16-bit thấp
        .slow_clk  (slow_clk)
    );

    // ------------------- Counter -------------------
    counter #(.WIDTH(WIDTH)) u_counter (
        .clk     (slow_clk),
        .rst_n   (rst_n),
        .PWM_EN  (en),
        .mode    (mode),
        .AAR     (period),
        .cnt_val (cnt_val)
    );

    // ------------------- Comparator -------------------
    comparator #(.WIDTH(WIDTH)) u_comparator (
        .CCR        (cnt_val),
        .CCR_COMPARE(duty),
        .period     (period),
        .enable     (en),
        .pwm_out    (PWM_OUT)
    );

endmodule
